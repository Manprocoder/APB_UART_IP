//==========================================================
//Project: Design APB-UART IP core
//File name: uvm_list.svh 
//Description: contains all UVM components
//==========================================================
//
//the line "import uvm_pkg::*" only impacts non-package files
//
`include "uvm_pkg.sv"
