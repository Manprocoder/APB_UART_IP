package parameter_pkg;
	parameter DW = 32;
	parameter APB_AW = 32;
	parameter OVERSAMPLE = 16;
endpackage

